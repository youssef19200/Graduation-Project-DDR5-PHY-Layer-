/**********************************************************************************
** Graduation project_S26
** Author: Ahmed Mohamed Zakaria
**
** Module Name: ddr5_phy_crc
** Description: this file contains the CRC Generation RTL (top module of the devices (X4, X8, X16))
**
*********************************************************************************/

module ddr5_phy_crc_gen 
    # (parameter pDRAM_SIZE = 4 )  // parameter indicate the device size (X4, X8, X16)
(
    // input signals //
	input 					clk_i ,         // clock signal
	input 					rst_n_i ,         // active low asynchronous reset
	input 					crc_en_i ,      // enable signal from write data block 
  	input  [2*pDRAM_SIZE-1: 0]	 crc_in_data_i , // input data bus from write data block that required crc code 
  
    // output signals //
  	output  [2*pDRAM_SIZE-1: 0]	 crc_code_o       // output crc bits 
);


    // duplicating crc block according to the device size
    genvar i ;

    generate
        for ( i=0 ; i< 2*pDRAM_SIZE ; i = i+8 )
	    begin
        ddr5_phy_crc_x4 crc_x4_U (
            .clk_i(clk_i),
            .rst_n_i(rst_n_i),
            .crc_en_i(crc_en_i),
            .crc_in_data_i (crc_in_data_i[i+7 : i]),
            .crc_code_o(crc_code_o[i+7 : i])
        );
	    end
  endgenerate

endmodule